`ifndef PP_CONSTANTS
`define PP_CONSTANTS
parameter NUM_SIZE=32;
parameter CMD_SIZE_LOG2=3;
`endif
