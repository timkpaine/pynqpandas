parameter NOOP=4'b0000;
parameter ADD=4'b0001;
