`ifndef DEF
`define DEF
parameter NOOP=4'b0000;
parameter ADD=4'b0001;
parameter NUM_SIZE=32;
parameter CMD_SIZE_LOG2=2;
`endif