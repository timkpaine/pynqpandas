`ifndef PP_DEF
`define PP_DEF
parameter NOOP=4'b0000;
parameter ADD=4'b0001;
parameter NUM_SIZE=32;
parameter CMD_SIZE_LOG2=3;
`endif