`ifndef DEF
`define DEF
parameter NOOP=4'b0000;
parameter ADD=4'b0001;
parameter NUM=31;
parameter CMD=3;
`endif