`ifndef PP_CONSTANTS
`define PP_CONSTANTS

`ifdef CC_MODELSIM
parameter NUM_SIZE=32;
parameter CMD_SIZE_LOG2=3;
`endif

`endif
