parameter NOOP=4'b0000;
